//----------------------------------------------------------------------------
//
//----------------------------------------------------------------------------
`timescale 1 ns / 100 ps

module system_tb;

//----------------------------------------------------------------------------
// Parameter (may differ for physical synthesis)
//----------------------------------------------------------------------------
parameter tck              = 10;       // clock period in ns
parameter uart_baud_rate   = 1152000;  // uart baud rate for simulation 

parameter clk_freq = 1000000000 / tck; // Frequenzy in HZ
//----------------------------------------------------------------------------
//
//----------------------------------------------------------------------------
reg        clk;
reg        rst;
//reg     [7:0]gpio0_io;     

/*wire       led;*/

//----------------------------------------------------------------------------
// UART STUFF (testbench uart, simulating a comm. partner)
//----------------------------------------------------------------------------
wire         uart_rxd;
wire         uart_txd;
wire	 [7:0]gpio_io;
reg     [7:0]gpio_dir;
reg     [7:0]data;


   genvar    i;
   generate 
      for (i=0;i<8;i=i+1)  begin: gpio_tris
	 assign gpio_io[i] = ~(gpio_dir[i]) ? data[i] : 1'bz;

	 end
   endgenerate

//----------------------------------------------------------------------------
// Device Under Test 
//----------------------------------------------------------------------------
system #(
	.clk_freq(           clk_freq         ),
	.uart_baud_rate(     uart_baud_rate   )
) dut  (
	.clk(          clk    ),
	// Debug
	.rst(          rst    ),
	/*.led(          led    ),*/
	// Uart
	.gpio0_io( gpio_io ),
	.uart_rxd(  uart_rxd  ),
	.uart_txd(  uart_txd  )
);


/* Clocking device */
initial         clk <= 0;
always #(tck/2) clk <= ~clk;

/* Simulation setup */
initial begin

        

	$dumpfile("system_tb.vcd");
	//$monitor("%b,%b,%b,%b",clk,rst,uart_txd,uart_rxd);
	$dumpvars(-1, dut);
	//$dumpvars(-1,clk,rst,uart_txd);
	// reset
	#0  rst <= 0;
	#100  rst <= 1;


	

	
	 

	#(tck*100000) $finish;
end



endmodule
